library verilog;
use verilog.vl_types.all;
entity MUX2to1TB is
end MUX2to1TB;
