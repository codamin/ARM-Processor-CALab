`timescale 1ns/1ns
module EXEStageTB();
  
endmodule
