library verilog;
use verilog.vl_types.all;
entity DataMemoryTB is
end DataMemoryTB;
