library verilog;
use verilog.vl_types.all;
entity InstructionMemoryTB is
end InstructionMemoryTB;
