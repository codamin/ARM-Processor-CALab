`timescale 1ns/1ns
module PCTB();
  
endmodule
