library verilog;
use verilog.vl_types.all;
entity PCTB is
end PCTB;
